//Same as q5a, but Mealy implementation
module top_module (
    input clk,
    input areset,
    input x,
    output z
); 
    parameter [1:0] A = 2'b01, B = 2'b10;
	reg [1:0] state, next;
	always @(*) begin
		case (state) 
			A : begin
				if (x) begin
					next = B;
					z =1;
				end
				else begin
					next = A;
					z = 0;
				end
			end
			B : begin
				next = B;
                z = (x) ? 1'b0 : 1'b1;
			end
		endcase
	end
    always @(posedge clk or posedge areset) begin
		if (areset) state <= A;
		else state <= next;
	end

endmodule
